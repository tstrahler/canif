library ieee;
use ieee.std_logic_1164.all;

entity top_tb is
end entity;

architecture top_tb_rtl of top_tb is

begin


end architecture;
